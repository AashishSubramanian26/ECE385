module datapath (	
                    input logic  LD_MAR, LD_MDR, LD_IR, LD_BEN, LD_CC, LD_REG, LD_PC, LD_LED, Clk, Reset, Run, Continue,
                    input logic  GatePC, GateMDR, GateALU, GateMARMUX,
                    input logic  SR2MUX, ADDR1MUX, MARMUX,
                    input logic  BEN, MIO_EN, DRMUX, SR1MUX,
                    input logic  [1:0] PCMUX, ADDR2MUX, ALUK,
                    input logic  [15:0] MDR_In,
					output logic [15:0]	MAR, MDR, IR //outputs
				);
				
	logic 	[15:0] 	BUS,
					IR_Reg_Out,
					MDR_Reg_Out,
					MAR_Out_Reg, 
					PC_Reg_Out, 
					MDR_MUX,
					PCMUX_Out;

	BusMux Tri_State_Buff(
					.S({GateMDR, GateALU, GatePC, GateMARMUX}), 
					.MARMUX(16'hxxxx), 
					.PC(PC_Reg_Out), 
					.ALU(16'hxxxx), 
					.MDR(MDR_Reg_Out), 
					.BUS(BUS)
					);

	Reg_16  MDR_Reg(
				.Clk(Clk),
				.Reset(Reset), 
				.Load(LD_MDR), 
				.D(MDR_MUX), 
				.Out(MDR_Reg_Out)
				);

	Reg_16  IR_Reg(
				.Clk(Clk),
				.Reset(Reset),	 
				.Load(LD_IR), 
				.D(BUS), 
				.Out(IR_Reg_Out)
				);

	Reg_16  PC_Reg(
				.Clk(Clk),
				.Reset(Reset),	 
				.Load(LD_PC), 
				.D(PCMUX_Out), 
				.Out(PC_Reg_Out)
				);

	Reg_16  MAR_Reg(
		.Clk(Clk),
		.Reset(Reset),	 
		.Load(LD_MAR), 
		.D(BUS), 
		.Out(MAR_Out_Reg)
		);

	TwoInputMux MDRMult (
				.S(MIO_EN), 
				.D1(BUS), 
				.D2(MDR_In), 
				.Out_Mux(MDR_MUX)
				);
	
	
	ThreeInputMux PCMult(
					.S(PCMUX), 
					.D3(PC_Reg_Out + 1'b1), 
					.D1(BUS), 
					.D2(16'hxxxx),
					.OUT(PCMUX_Out)
					);

	always_comb begin
		MDR_out = MDR_Reg_Out;
		MAR_out = MAR_Out_Reg;
		IR_out = IR_Reg_Out;
		PC_out = PC_Reg_Out;
	end 
endmodule 