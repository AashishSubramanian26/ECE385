module register_unit (input  logic Clk, A_In, B_In, Ld_A, Ld_B, 
                            Shift_En, Reset, ClearXA,
                      input  logic [7:0]  D_A, D_B, 
                      output logic A_out, B_out, 
                      output logic [7:0]  A,
                      output logic [7:0]  B);


    reg_8  reg_A (.Clk(Clk), .Reset(Reset | ClearXA), .Shift_In(A_In), .Load(Ld_A), .Shift_En(Shift_En),
	               .D(D_A), .Shift_Out(A_out), .Data_Out(A));
    reg_8  reg_B (.Clk(Clk), .Reset(1'b0), .Shift_In(B_In), .Load(Reset), .Shift_En(Shift_En),
	               .D(D_B), .Shift_Out(B_out), .Data_Out(B));

endmodule