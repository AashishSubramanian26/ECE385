module testbench();

timeunit 10ns;

timeprecision 1ns;